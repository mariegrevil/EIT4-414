library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
--use ieee.std_logic_unsigned.all;

entity TestBench is

	--port(

		--);
end TestBench;

architecture rtl of TestBench is

begin

end rtl;