library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ProgramCode is
    port (TinyClock  		: in std_logic;
          DataBusProgram	: out std_logic_vector(31 downto 0); -- Data on the chosen addres
		  AddrBusProgram	: in std_logic_vector(7 downto 0); -- The addres that the CU wants to load
		  ClockCycle 		: in std_logic_vector(2 downto 0) -- Counts rising edges in tinyclock per hugeclock
		  ); 
		  
end  ProgramCode;

architecture rtl of Programcode is

    type ProMem_type is array (255 downto 0) of std_logic_vector (31 downto 0); -- Declare a data type. here an array with 255 locations of 32 bits
    signal ProMem: ProMem_type := (others => x"00000000"); -- A signal of type "ProMem_type". All values are preconfigured to 0
	
begin
-- ActionJackson-værdier:
-- 17 er plus+facit
-- 9 er minus+facit
-- 5 er gange+facit
-- 3 er divider+facit

ProMem(0) <= "00101000001111000000000000000001"; -- SET 30 REG 0
ProMem(1) <= "00101000001101100000000000000001"; -- SET 27 REG 0
-- MARK start at ProMem(2)
ProMem(2) <= "01001000000000011111100000100011"; -- BNEQ 31 17
ProMem(3) <= "10110000000000010000000000010111"; -- GOTO plus
ProMem(4) <= "01001000000000011111100000010011"; -- BNEQ 31 9
ProMem(5) <= "10110000000000010000000000011101"; -- GOTO minus
ProMem(6) <= "01001000000000011111100000001011"; -- BNEQ 31 5
ProMem(7) <= "10110000000000010000000000100011"; -- GOTO gange
ProMem(8) <= "01001000000000011111100000000111"; -- BNEQ 31 3
ProMem(9) <= "10110000000000010000000000101001"; -- GOTO divider
ProMem(10) <= "10110000000000010000000000000101"; -- GOTO start
-- MARK plus at ProMem(11)
ProMem(11) <= "01010000001111001110000000111010"; -- ADD 30 REG 28 29 REG
ProMem(12) <= "11111000001101100000000000000001"; -- TBR 27 REG 
ProMem(13) <= "10110000000000010000000000101111"; -- GOTO clear
-- MARK minus at ProMem(14)
ProMem(14) <= "01100000001111001110000000111010"; -- SUB 30 REG 28 29 REG
ProMem(15) <= "11111000001101100000000000000001"; -- TBR 27 REG 
ProMem(16) <= "10110000000000010000000000101111"; -- GOTO clear
-- MARK gange at ProMem(17)
ProMem(17) <= "01110000001111001110000000111010"; -- MULT 30 REG 28 29 REG
ProMem(18) <= "11111000001101100000000000000001"; -- TBR 27 REG 
ProMem(19) <= "10110000000000010000000000101111"; -- GOTO clear
-- MARK divider at ProMem(20)
ProMem(20) <= "01111000001111001110000000111010"; -- DIV 30 REG 28 29 REG
ProMem(21) <= "11111000001101100000000000000001"; -- TBR 27 REG 
ProMem(22) <= "10110000000000010000000000101111"; -- GOTO clear
-- MARK clear at ProMem(23)
ProMem(23) <= "01000000000000011111100001000001"; -- BEQ 31 32
ProMem(24) <= "10111000000000010000000000000011"; -- JMPX 1
ProMem(25) <= "00101000001111000000000000000001"; -- SET 30 REG 0
ProMem(26) <= "00101000001101100000000000000001"; -- SET 27 REG 0
ProMem(27) <= "10110000000000010000000000000101"; -- GOTO start

-- Interrupt 1 "rest"
ProMem(28) <= "00101000000000000000000000000001"; -- SET 0 REG 0
ProMem(29) <= "00101000000000100000000000000001"; -- SET 1 REG 0
ProMem(30) <= "00101000000001000000000000000001"; -- SET 2 REG 0
ProMem(31) <= "00101000000001100000000000000001"; -- SET 3 REG 0
ProMem(32) <= "00101000000010000000000000000001"; -- SET 4 REG 0
ProMem(33) <= "00101000000010100000000000000001"; -- SET 5 REG 0
ProMem(34) <= "00101000000011000000000000000001"; -- SET 6 REG 0
ProMem(35) <= "00101000000011100000000000000001"; -- SET 7 REG 0
ProMem(36) <= "00101000000100000000000000000001"; -- SET 8 REG 0
ProMem(37) <= "00101000000100100000000000000001"; -- SET 9 REG 0
ProMem(38) <= "00101000000101000000000000000001"; -- SET 10 REG 0
ProMem(39) <= "00101000000101100000000000000001"; -- SET 11 REG 0
ProMem(40) <= "00101000000110000000000000000001"; -- SET 12 REG 0
ProMem(41) <= "00101000000110100000000000000001"; -- SET 13 REG 0
ProMem(42) <= "00101000000111000000000000000001"; -- SET 14 REG 0
ProMem(43) <= "00101000000111100000000000000001"; -- SET 15 REG 0
ProMem(44) <= "00101000001000000000000000000001"; -- SET 16 REG 0
ProMem(45) <= "00101000001000100000000000000001"; -- SET 17 REG 0
ProMem(46) <= "00101000001001000000000000000001"; -- SET 18 REG 0
ProMem(47) <= "00101000001001100000000000000001"; -- SET 19 REG 0
ProMem(48) <= "00101000001010000000000000000001"; -- SET 20 REG 0
ProMem(49) <= "00101000001010100000000000000001"; -- SET 21 REG 0
ProMem(50) <= "00101000001011000000000000000001"; -- SET 22 REG 0
ProMem(51) <= "00101000001011100000000000000001"; -- SET 23 REG 0
ProMem(52) <= "00101000001100000000000000000001"; -- SET 24 REG 0
ProMem(53) <= "00101000001100100000000000000001"; -- SET 25 REG 0
ProMem(54) <= "00101000001101000000000000000001"; -- SET 26 REG 0
ProMem(55) <= "00101000001101100000000000000001"; -- SET 27 REG 0
ProMem(56) <= "00101000001110000000000000000001"; -- SET 28 REG 0
ProMem(57) <= "00101000001110100000000000000001"; -- SET 29 REG 0
ProMem(58) <= "00101000001110000000000000000001"; -- SET 28 REG 0
ProMem(59) <= "00101000001110100000000000000001"; -- SET 29 REG 0
ProMem(60) <= "00101000001111000000000000000001"; -- SET 30 REG 0
ProMem(61) <= "00101000001111100000000000000001"; -- SET 31 REG 0
ProMem(62) <= "10110000000000010000000000000101"; -- GOTO start

			
process (TinyClock)
    begin
	if Clockcycle = "001" then 
        if rising_edge(TinyClock) then
            DataBusProgram <= ProMem(conv_integer(AddrBusProgram));  --Put the location pointet to by the "AddrBusProgram" on to "DataBusProgram"
            
        end if;
	end if;
    end process;

end rtl;
